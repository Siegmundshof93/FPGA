module div_clk
(
input clk,


output reg d_clk
);

 reg [23:0] count = 24'b0;
 reg [23:0] COUNT_MAX = 24'd12000000;

always @ (posedge clk)
begin
 if(count == COUNT_MAX)
    begin
      count <= 24'b0;
      d_clk <= ~d_clk;
    end
    else
      begin
    count <= count + 1;
      end
end

endmodule
